*** SPICE deck for cell OR{sch} from library term_project
*** Created on Cmt Ara 24, 2022 15:48:05
*** Last revised on Sal Ara 27, 2022 14:44:10
*** Written on Çar Ara 28, 2022 13:43:14 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT term_project__NOR__FOR_OR_ FROM CELL NOR_(FOR_OR){sch}
.SUBCKT term_project__NOR__FOR_OR_ A AnorB B
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 AnorB A gnd gnd NMOS L=0.36U W=0.9U
Mnmos@1 AnorB B gnd gnd NMOS L=0.36U W=0.9U
Mpmos@0 AnorB B net@19 vdd PMOS L=0.36U W=3.6U
Mpmos@1 net@19 A vdd vdd PMOS L=0.36U W=3.6U
.ENDS term_project__NOR__FOR_OR_

*** SUBCIRCUIT term_project__inverter FROM CELL inverter{sch}
.SUBCKT term_project__inverter A notA
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 notA A gnd gnd NMOS L=0.36U W=0.9U
Mpmos@0 notA A vdd vdd PMOS L=0.36U W=1.8U
.ENDS term_project__inverter

.global gnd vdd

*** TOP LEVEL CELL: OR{sch}
XNOR@2 A net@0 B term_project__NOR__FOR_OR_
Xinverter@0 net@0 AorB term_project__inverter

* Spice Code nodes in cell cell 'OR{sch}'
vdd vdd 0 dc 5
va A 0 DC 0 pulse 0 5 1n 1n 1n 10m 20m
vb B 0 DC 0 pulse 0 5 1n 1n 1n 5m 10m
.tran 0 20m
.include /Applications/electric_vlsi/process/C5_models.txt
.END
