*** SPICE deck for cell XOR{sch} from library term_project
*** Created on Pzt Ara 26, 2022 08:55:50
*** Last revised on Sal Ara 27, 2022 14:45:30
*** Written on Sal Ara 27, 2022 14:45:36 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

.global gnd vdd

*** TOP LEVEL CELL: XOR{sch}
Mnmos@0 net@1 B gnd gnd N L=0.36U W=0.9U
Mnmos@1 net@1 A AxorB gnd N L=0.36U W=0.9U
Mnmos@2 B net@13 AxorB gnd N L=0.36U W=0.9U
Mnmos@3 net@13 A gnd gnd N L=0.36U W=0.9U
Mpmos@0 vdd B net@1 vdd P L=0.36U W=1.8U
Mpmos@1 net@1 net@13 AxorB vdd P L=0.36U W=1.8U
Mpmos@2 B A AxorB vdd P L=0.36U W=1.8U
Mpmos@3 vdd A net@13 vdd P L=0.36U W=1.8U

* Spice Code nodes in cell cell 'XOR{sch}'
vdd vdd 0 dc 5
va A 0 DC 0 pulse 0 5 1n 1n 1n 10m 20m
vb B 0 DC 0 pulse 0 5 1n 1n 1n 5m 10m
.tran 0 20m
.include /Applications/electric_vlsi/process/C5_models.txt
.END
