*** SPICE deck for cell 3NAND{sch} from library term_project
*** Created on Per Eki 06, 2022 17:52:59
*** Last revised on Per Ara 29, 2022 15:23:26
*** Written on Per Ara 29, 2022 15:36:08 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

.global gnd vdd

*** TOP LEVEL CELL: 3NAND{sch}
Mnmos@1 ABC A net@15 gnd NMOS L=0.36U W=1.8U
Mnmos@2 net@15 B net@33 gnd NMOS L=0.36U W=1.8U
Mnmos@3 net@33 C gnd gnd NMOS L=0.36U W=1.8U
Mpmos@0 ABC A vdd vdd PMOS L=0.36U W=1.8U
Mpmos@1 ABC B vdd vdd PMOS L=0.36U W=1.8U
Mpmos@2 ABC C vdd vdd PMOS L=0.36U W=1.8U

* Spice Code nodes in cell cell '3NAND{sch}'
vdd vdd 0 dc 5
va A 0 DC 0 pulse 0 5 1n 1n 1n 20m 40m
vb B 0 DC 0 pulse 0 5 1n 1n 1n 10m 20m
vc C 0 DC 0 pulse 0 5 1n 1n 1n 5m 10m
.tran 0 40m
.include /Applications/electric_vlsi/process/C5_models.txt
.END
