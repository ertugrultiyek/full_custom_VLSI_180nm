*** SPICE deck for cell ALU_Mid_Bits{sch} from library term_project_backup_00
*** Created on Cum Ara 30, 2022 04:05:23
*** Last revised on Cum Ara 30, 2022 18:29:11
*** Written on Per Oca 05, 2023 14:15:23 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT term_project_backup_00__3NAND FROM CELL 3NAND{sch}
.SUBCKT term_project_backup_00__3NAND A ABC_ B C
** GLOBAL gnd
** GLOBAL vdd
Mnmos@1 ABC_ A net@15 gnd NMOS L=0.36U W=1.8U
Mnmos@2 net@15 B net@33 gnd NMOS L=0.36U W=1.8U
Mnmos@3 net@33 C gnd gnd NMOS L=0.36U W=1.8U
Mpmos@0 ABC_ A vdd vdd PMOS L=0.36U W=1.8U
Mpmos@1 ABC_ B vdd vdd PMOS L=0.36U W=1.8U
Mpmos@2 ABC_ C vdd vdd PMOS L=0.36U W=1.8U
.ENDS term_project_backup_00__3NAND

*** SUBCIRCUIT term_project_backup_00__inverter FROM CELL inverter{sch}
.SUBCKT term_project_backup_00__inverter A notA
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 notA A gnd gnd NMOS L=0.36U W=0.9U
Mpmos@0 notA A vdd vdd PMOS L=0.36U W=1.8U
.ENDS term_project_backup_00__inverter

*** SUBCIRCUIT term_project_backup_00__3NAND/AND FROM CELL 3NAND/AND{sch}
.SUBCKT term_project_backup_00__3NAND/AND A ABC ABC_ B C
** GLOBAL gnd
** GLOBAL vdd
X_3NAND@1 A ABC_ B C term_project_backup_00__3NAND
Xinverter@0 ABC_ ABC term_project_backup_00__inverter
.ENDS term_project_backup_00__3NAND/AND

*** SUBCIRCUIT term_project_backup_00__NAND FROM CELL NAND{sch}
.SUBCKT term_project_backup_00__NAND A AnandB B
** GLOBAL gnd
** GLOBAL vdd
Mnmos@1 AnandB A net@15 gnd NMOS L=0.36U W=1.8U
Mnmos@2 net@15 B gnd gnd NMOS L=0.36U W=1.8U
Mpmos@0 AnandB A vdd vdd PMOS L=0.36U W=1.8U
Mpmos@1 AnandB B vdd vdd PMOS L=0.36U W=1.8U
.ENDS term_project_backup_00__NAND

*** SUBCIRCUIT term_project_backup_00__AND FROM CELL AND{sch}
.SUBCKT term_project_backup_00__AND A AandB B
** GLOBAL gnd
** GLOBAL vdd
XNAND@0 A net@2 B term_project_backup_00__NAND
Xinverter@0 net@2 AandB term_project_backup_00__inverter
.ENDS term_project_backup_00__AND

*** SUBCIRCUIT term_project_backup_00__Multiplexer FROM CELL Multiplexer{sch}
.SUBCKT term_project_backup_00__Multiplexer A B F notS S
** GLOBAL gnd
** GLOBAL vdd
Mnmos@7 F notS B gnd N L=0.36U W=1.8U
Mnmos@8 F S A gnd N L=0.36U W=1.8U
Mpmos@7 F S B vdd P L=0.36U W=1.8U
Mpmos@8 F notS A vdd P L=0.36U W=1.8U
.ENDS term_project_backup_00__Multiplexer

*** SUBCIRCUIT term_project_backup_00__NAND/AND FROM CELL NAND/AND{sch}
.SUBCKT term_project_backup_00__NAND/AND A AandB AnandB B
** GLOBAL gnd
** GLOBAL vdd
XNAND@0 A AnandB B term_project_backup_00__NAND
Xinverter@0 AnandB AandB term_project_backup_00__inverter
.ENDS term_project_backup_00__NAND/AND

*** SUBCIRCUIT term_project_backup_00__XOR FROM CELL XOR{sch}
.SUBCKT term_project_backup_00__XOR A AxorB B
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 net@1 B gnd gnd N L=0.36U W=0.9U
Mnmos@1 net@1 A AxorB gnd N L=0.36U W=0.9U
Mnmos@2 B net@13 AxorB gnd N L=0.36U W=0.9U
Mnmos@3 net@13 A gnd gnd N L=0.36U W=0.9U
Mpmos@0 vdd B net@1 vdd P L=0.36U W=1.8U
Mpmos@1 net@1 net@13 AxorB vdd P L=0.36U W=1.8U
Mpmos@2 B A AxorB vdd P L=0.36U W=1.8U
Mpmos@3 vdd A net@13 vdd P L=0.36U W=1.8U
.ENDS term_project_backup_00__XOR

*** SUBCIRCUIT term_project_backup_00__Half_Adder FROM CELL Half_Adder{sch}
.SUBCKT term_project_backup_00__Half_Adder A A+B B Cout
** GLOBAL gnd
** GLOBAL vdd
XAND@0 A Cout B term_project_backup_00__AND
XXOR@2 B A+B A term_project_backup_00__XOR
.ENDS term_project_backup_00__Half_Adder

*** SUBCIRCUIT term_project_backup_00__NOR__FOR_OR_ FROM CELL NOR_(FOR_OR){sch}
.SUBCKT term_project_backup_00__NOR__FOR_OR_ A AnorB B
** GLOBAL gnd
** GLOBAL vdd
Mnmos@0 AnorB A gnd gnd NMOS L=0.36U W=0.9U
Mnmos@1 AnorB B gnd gnd NMOS L=0.36U W=0.9U
Mpmos@0 AnorB B net@19 vdd PMOS L=0.36U W=3.6U
Mpmos@1 net@19 A vdd vdd PMOS L=0.36U W=3.6U
.ENDS term_project_backup_00__NOR__FOR_OR_

*** SUBCIRCUIT term_project_backup_00__OR FROM CELL OR{sch}
.SUBCKT term_project_backup_00__OR A AorB B
** GLOBAL gnd
** GLOBAL vdd
XNOR@2 A net@0 B term_project_backup_00__NOR__FOR_OR_
Xinverter@0 net@0 AorB term_project_backup_00__inverter
.ENDS term_project_backup_00__OR

*** SUBCIRCUIT term_project_backup_00__Full_Adder FROM CELL Full_Adder{sch}
.SUBCKT term_project_backup_00__Full_Adder A A+B B Cin Cout
** GLOBAL gnd
** GLOBAL vdd
XHalf_Add@0 A net@0 B net@12 term_project_backup_00__Half_Adder
XHalf_Add@1 net@0 A+B Cin net@17 term_project_backup_00__Half_Adder
XOR@1 net@12 Cout net@17 term_project_backup_00__OR
.ENDS term_project_backup_00__Full_Adder

*** SUBCIRCUIT term_project_backup_00__adder_subtractor FROM CELL adder_subtractor{sch}
.SUBCKT term_project_backup_00__adder_subtractor A B C/B_in C/B_out operator Result
** GLOBAL gnd
** GLOBAL vdd
XFull_Add@0 A Result net@0 C/B_in C/B_out term_project_backup_00__Full_Adder
XXOR@0 operator net@0 B term_project_backup_00__XOR
.ENDS term_project_backup_00__adder_subtractor

*** SUBCIRCUIT term_project_backup_00__AU_mid FROM CELL AU_mid{sch}
.SUBCKT term_project_backup_00__AU_mid A B C/B_out Cin Cout_inp notCin notS0 notS2 result S1 S2
** GLOBAL gnd
** GLOBAL vdd
X_3NAND/AN@0 notCin net@125 net@124 notS0 notS2 term_project_backup_00__3NAND/AND
X_3NAND@0 notS2 net@44 notS0 Cin term_project_backup_00__3NAND
XMultiple@0 gnd B net@5 net@137 net@139 term_project_backup_00__Multiplexer
XMultiple@1 gnd Cout_inp net@55 net@124 net@125 term_project_backup_00__Multiplexer
XNAND/AND@0 net@44 net@139 net@137 net@45 term_project_backup_00__NAND/AND
XNAND@0 S1 net@45 S2 term_project_backup_00__NAND
Xadder_su@0 A net@5 net@55 C/B_out S2 result term_project_backup_00__adder_subtractor
.ENDS term_project_backup_00__AU_mid

*** SUBCIRCUIT term_project_backup_00__NOR/OR FROM CELL NOR/OR{sch}
.SUBCKT term_project_backup_00__NOR/OR A AnorB AorB B
** GLOBAL gnd
** GLOBAL vdd
XNOR@2 A AnorB B term_project_backup_00__NOR__FOR_OR_
Xinverter@0 AnorB AorB term_project_backup_00__inverter
.ENDS term_project_backup_00__NOR/OR

*** SUBCIRCUIT term_project_backup_00__D_LATCH FROM CELL D_LATCH{sch}
.SUBCKT term_project_backup_00__D_LATCH clk D notQ Q
** GLOBAL gnd
** GLOBAL vdd
XMultiple@0 D Q net@1 net@14 clk term_project_backup_00__Multiplexer
Xinverter@0 net@1 notQ term_project_backup_00__inverter
Xinverter@1 notQ Q term_project_backup_00__inverter
Xinverter@2 clk net@14 term_project_backup_00__inverter
.ENDS term_project_backup_00__D_LATCH

*** SUBCIRCUIT term_project_backup_00__D_FF FROM CELL D_FF{sch}
.SUBCKT term_project_backup_00__D_FF clk D notQ Q
** GLOBAL gnd
** GLOBAL vdd
XD_LATCH@0 clk D D_LATCH@0_notQ net@0 term_project_backup_00__D_LATCH
XD_LATCH@1 net@1 net@0 notQ Q term_project_backup_00__D_LATCH
Xinverter@0 clk net@1 term_project_backup_00__inverter
.ENDS term_project_backup_00__D_FF

*** SUBCIRCUIT term_project_backup_00__Shift_Register FROM CELL Shift_Register{sch}
.SUBCKT term_project_backup_00__Shift_Register clk Dir F L notDir R
** GLOBAL gnd
** GLOBAL vdd
XD_FF@0 clk net@8 D_FF@0_notQ F term_project_backup_00__D_FF
XMultiple@0 R L net@8 notDir Dir term_project_backup_00__Multiplexer
.ENDS term_project_backup_00__Shift_Register

.global gnd vdd

*** TOP LEVEL CELL: ALU_Mid_Bits{sch}
X_3NAND/AN@0 S0 net@89 net@92 S2 S1 term_project_backup_00__3NAND/AND
XAND@0 net@14 net@9 B term_project_backup_00__AND
XAU_mid@0 net@14 B C/B_out Cin C/B_in notCin notS0 notS2 net@58 S1 S2 term_project_backup_00__AU_mid
XMultiple@0 net@14 net@2 net@35 Cin notCin term_project_backup_00__Multiplexer
XMultiple@1 net@9 net@10 net@38 Cin notCin term_project_backup_00__Multiplexer
XMultiple@2 net@55 net@58 net@48 net@92 net@89 term_project_backup_00__Multiplexer
XMultiple@3 net@35 net@38 net@43 S0 notS0 term_project_backup_00__Multiplexer
XMultiple@4 net@43 net@48 F net@52 net@53 term_project_backup_00__Multiplexer
XNOR/OR@0 S1 net@53 net@52 S2 term_project_backup_00__NOR/OR
XOR@0 net@14 net@10 B term_project_backup_00__OR
XShift_Re@0 clk Cin net@55 L notCin R term_project_backup_00__Shift_Register
Xinverter@0 A net@2 term_project_backup_00__inverter
Xinverter@1 net@2 net@14 term_project_backup_00__inverter

* Spice Code nodes in cell cell 'ALU_Mid_Bits{sch}'
vdd vdd 0 dc 5
vs2 S2 0 DC 0 pulse 5 0 1n 1n 1n 256m 512m
vns2 notS2 0 DC 0 pulse 0 5 1n 1n 1n 256m 512m
vs1 S1 0 DC 0 pulse 5 0 1n 1n 1n 128m 256m
vns1 notS1 0 DC 0 pulse 0 5 1n 1n 1n 128m 256m
vs0 S0 0 DC 0 pulse 5 0 1n 1n 1n 64m 128m
vns0 notS0 0 DC 0 pulse 0 5 1n 1n 1n 64m 128m
vcin Cin 0 DC 0 pulse 5 0 1n 1n 1n 32m 64m
vncin notCin 0 DC 0 pulse 0 5 1n 1n 1n 32m 64m
vcb_in C/B_in 0 DC 0 pulse 5 0 1n 1n 1n 16m 32m
va A 0 DC 0 pulse 5 0 1n 1n 1n 8m 16m
vb B 0 DC 0 pulse 5 0 1n 1n 1n 4m 8m
vl L 0 DC 0 pulse 5 0 1n 1n 1n 2m 4m
vr R 0 DC 0 pulse 5 0 1n 1n 1n 1m 2m
vclk clk 0 DC 0 pulse 5 0 1n 1n 1n 0.4m 1m
.tran 0 512m
.include /Applications/electric_vlsi/process/C5_models.txt
.END
